// Verilog
// c1355
// Ninputs 41
// Noutputs 32
// NtotalGates 546
// AND2 40
// NAND2 416
// NOT1 40
// AND4 8
// OR4 2
// AND5 8
// BUFF1 32

module c1355 (N1,N8,N15,N22,N29,N36,N43,N50,N57,N64,
              N71,N78,N85,N92,N99,N106,N113,N120,N127,N134,
              N141,N148,N155,N162,N169,N176,N183,N190,N197,N204,
              N211,N218,N225,N226,N227,N228,N229,N230,N231,N232,
              N233,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,
              N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
              N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
              N1353,N1354,N1355);

input N1,N8,N15,N22,N29,N36,N43,N50,N57,N64,
      N71,N78,N85,N92,N99,N106,N113,N120,N127,N134,
      N141,N148,N155,N162,N169,N176,N183,N190,N197,N204,
      N211,N218,N225,N226,N227,N228,N229,N230,N231,N232,
      N233;

output N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,
       N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
       N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
       N1354,N1355;

wire N242,N245,N248,N251,N254,N257,N260,N263,N266,N269,
     N272,N275,N278,N281,N284,N287,N290,N293,N296,N299,
     N302,N305,N308,N311,N314,N317,N320,N323,N326,N329,
     N332,N335,N338,N341,N344,N347,N350,N353,N356,N359,
     N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
     N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
     N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,
     N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,
     N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,
     N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
     N422,N423,N424,N425,N426,N429,N432,N435,N438,N441,
     N444,N447,N450,N453,N456,N459,N462,N465,N468,N471,
     N474,N477,N480,N483,N486,N489,N492,N495,N498,N501,
     N504,N507,N510,N513,N516,N519,N522,N525,N528,N531,
     N534,N537,N540,N543,N546,N549,N552,N555,N558,N561,
     N564,N567,N570,N571,N572,N573,N574,N575,N576,N577,
     N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,
     N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
     N598,N599,N600,N601,N602,N607,N612,N617,N622,N627,
     N632,N637,N642,N645,N648,N651,N654,N657,N660,N663,
     N666,N669,N672,N675,N678,N681,N684,N687,N690,N691,
     N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,
     N702,N703,N704,N705,N706,N709,N712,N715,N718,N721,
     N724,N727,N730,N733,N736,N739,N742,N745,N748,N751,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N767,N768,N769,N770,N773,N776,N779,
     N782,N785,N788,N791,N794,N797,N800,N803,N806,N809,
     N812,N815,N818,N819,N820,N821,N822,N823,N824,N825,
     N826,N827,N828,N829,N830,N831,N832,N833,N834,N847,
     N860,N873,N886,N899,N912,N925,N938,N939,N940,N941,
     N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,
     N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,
     N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,
     N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
     N982,N983,N984,N985,N986,N991,N996,N1001,N1006,N1011,
     N1016,N1021,N1026,N1031,N1036,N1039,N1042,N1045,N1048,N1051,
     N1054,N1057,N1060,N1063,N1066,N1069,N1072,N1075,N1078,N1081,
     N1084,N1087,N1090,N1093,N1096,N1099,N1102,N1105,N1108,N1111,
     N1114,N1117,N1120,N1123,N1126,N1129,N1132,N1135,N1138,N1141,
     N1144,N1147,N1150,N1153,N1156,N1159,N1162,N1165,N1168,N1171,
     N1174,N1177,N1180,N1183,N1186,N1189,N1192,N1195,N1198,N1201,
     N1204,N1207,N1210,N1213,N1216,N1219,N1222,N1225,N1228,N1229,
     N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,
     N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
     N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,
     N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,
     N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,
     N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
     N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,
     N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,
     N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,
     N1320,N1321,N1322,N1323;

and AND2_1 (N242, N225, N233);
and AND2_2 (N245, N226, N233);
and AND2_3 (N248, N227, N233);
and AND2_4 (N251, N228, N233);
and AND2_5 (N254, N229, N233);
and AND2_6 (N257, N230, N233);
and AND2_7 (N260, N231, N233);
and AND2_8 (N263, N232, N233);
nand NAND2_9 (N266, N1, N8);
nand NAND2_10 (N269, N15, N22);
nand NAND2_11 (N272, N29, N36);
nand NAND2_12 (N275, N43, N50);
nand NAND2_13 (N278, N57, N64);
nand NAND2_14 (N281, N71, N78);
nand NAND2_15 (N284, N85, N92);
nand NAND2_16 (N287, N99, N106);
nand NAND2_17 (N290, N113, N120);
nand NAND2_18 (N293, N127, N134);
nand NAND2_19 (N296, N141, N148);
nand NAND2_20 (N299, N155, N162);
nand NAND2_21 (N302, N169, N176);
nand NAND2_22 (N305, N183, N190);
nand NAND2_23 (N308, N197, N204);
nand NAND2_24 (N311, N211, N218);
nand NAND2_25 (N314, N1, N29);
nand NAND2_26 (N317, N57, N85);
nand NAND2_27 (N320, N8, N36);
nand NAND2_28 (N323, N64, N92);
nand NAND2_29 (N326, N15, N43);
nand NAND2_30 (N329, N71, N99);
nand NAND2_31 (N332, N22, N50);
nand NAND2_32 (N335, N78, N106);
nand NAND2_33 (N338, N113, N141);
nand NAND2_34 (N341, N169, N197);
nand NAND2_35 (N344, N120, N148);
nand NAND2_36 (N347, N176, N204);
nand NAND2_37 (N350, N127, N155);
nand NAND2_38 (N353, N183, N211);
nand NAND2_39 (N356, N134, N162);
nand NAND2_40 (N359, N190, N218);
nand NAND2_41 (N362, N1, N266);
nand NAND2_42 (N363, N8, N266);
nand NAND2_43 (N364, N15, N269);
nand NAND2_44 (N365, N22, N269);
nand NAND2_45 (N366, N29, N272);
nand NAND2_46 (N367, N36, N272);
nand NAND2_47 (N368, N43, N275);
nand NAND2_48 (N369, N50, N275);
nand NAND2_49 (N370, N57, N278);
nand NAND2_50 (N371, N64, N278);
nand NAND2_51 (N372, N71, N281);
nand NAND2_52 (N373, N78, N281);
nand NAND2_53 (N374, N85, N284);
nand NAND2_54 (N375, N92, N284);
nand NAND2_55 (N376, N99, N287);
nand NAND2_56 (N377, N106, N287);
nand NAND2_57 (N378, N113, N290);
nand NAND2_58 (N379, N120, N290);
nand NAND2_59 (N380, N127, N293);
nand NAND2_60 (N381, N134, N293);
nand NAND2_61 (N382, N141, N296);
nand NAND2_62 (N383, N148, N296);
nand NAND2_63 (N384, N155, N299);
nand NAND2_64 (N385, N162, N299);
nand NAND2_65 (N386, N169, N302);
nand NAND2_66 (N387, N176, N302);
nand NAND2_67 (N388, N183, N305);
nand NAND2_68 (N389, N190, N305);
nand NAND2_69 (N390, N197, N308);
nand NAND2_70 (N391, N204, N308);
nand NAND2_71 (N392, N211, N311);
nand NAND2_72 (N393, N218, N311);
nand NAND2_73 (N394, N1, N314);
nand NAND2_74 (N395, N29, N314);
nand NAND2_75 (N396, N57, N317);
nand NAND2_76 (N397, N85, N317);
nand NAND2_77 (N398, N8, N320);
nand NAND2_78 (N399, N36, N320);
nand NAND2_79 (N400, N64, N323);
nand NAND2_80 (N401, N92, N323);
nand NAND2_81 (N402, N15, N326);
nand NAND2_82 (N403, N43, N326);
nand NAND2_83 (N404, N71, N329);
nand NAND2_84 (N405, N99, N329);
nand NAND2_85 (N406, N22, N332);
nand NAND2_86 (N407, N50, N332);
nand NAND2_87 (N408, N78, N335);
nand NAND2_88 (N409, N106, N335);
nand NAND2_89 (N410, N113, N338);
nand NAND2_90 (N411, N141, N338);
nand NAND2_91 (N412, N169, N341);
nand NAND2_92 (N413, N197, N341);
nand NAND2_93 (N414, N120, N344);
nand NAND2_94 (N415, N148, N344);
nand NAND2_95 (N416, N176, N347);
nand NAND2_96 (N417, N204, N347);
nand NAND2_97 (N418, N127, N350);
nand NAND2_98 (N419, N155, N350);
nand NAND2_99 (N420, N183, N353);
nand NAND2_100 (N421, N211, N353);
nand NAND2_101 (N422, N134, N356);
nand NAND2_102 (N423, N162, N356);
nand NAND2_103 (N424, N190, N359);
nand NAND2_104 (N425, N218, N359);
nand NAND2_105 (N426, N362, N363);
nand NAND2_106 (N429, N364, N365);
nand NAND2_107 (N432, N366, N367);
nand NAND2_108 (N435, N368, N369);
nand NAND2_109 (N438, N370, N371);
nand NAND2_110 (N441, N372, N373);
nand NAND2_111 (N444, N374, N375);
nand NAND2_112 (N447, N376, N377);
nand NAND2_113 (N450, N378, N379);
nand NAND2_114 (N453, N380, N381);
nand NAND2_115 (N456, N382, N383);
nand NAND2_116 (N459, N384, N385);
nand NAND2_117 (N462, N386, N387);
nand NAND2_118 (N465, N388, N389);
nand NAND2_119 (N468, N390, N391);
nand NAND2_120 (N471, N392, N393);
nand NAND2_121 (N474, N394, N395);
nand NAND2_122 (N477, N396, N397);
nand NAND2_123 (N480, N398, N399);
nand NAND2_124 (N483, N400, N401);
nand NAND2_125 (N486, N402, N403);
nand NAND2_126 (N489, N404, N405);
nand NAND2_127 (N492, N406, N407);
nand NAND2_128 (N495, N408, N409);
nand NAND2_129 (N498, N410, N411);
nand NAND2_130 (N501, N412, N413);
nand NAND2_131 (N504, N414, N415);
nand NAND2_132 (N507, N416, N417);
nand NAND2_133 (N510, N418, N419);
nand NAND2_134 (N513, N420, N421);
nand NAND2_135 (N516, N422, N423);
nand NAND2_136 (N519, N424, N425);
nand NAND2_137 (N522, N426, N429);
nand NAND2_138 (N525, N432, N435);
nand NAND2_139 (N528, N438, N441);
nand NAND2_140 (N531, N444, N447);
nand NAND2_141 (N534, N450, N453);
nand NAND2_142 (N537, N456, N459);
nand NAND2_143 (N540, N462, N465);
nand NAND2_144 (N543, N468, N471);
nand NAND2_145 (N546, N474, N477);
nand NAND2_146 (N549, N480, N483);
nand NAND2_147 (N552, N486, N489);
nand NAND2_148 (N555, N492, N495);
nand NAND2_149 (N558, N498, N501);
nand NAND2_150 (N561, N504, N507);
nand NAND2_151 (N564, N510, N513);
nand NAND2_152 (N567, N516, N519);
nand NAND2_153 (N570, N426, N522);
nand NAND2_154 (N571, N429, N522);
nand NAND2_155 (N572, N432, N525);
nand NAND2_156 (N573, N435, N525);
nand NAND2_157 (N574, N438, N528);
nand NAND2_158 (N575, N441, N528);
nand NAND2_159 (N576, N444, N531);
nand NAND2_160 (N577, N447, N531);
nand NAND2_161 (N578, N450, N534);
nand NAND2_162 (N579, N453, N534);
nand NAND2_163 (N580, N456, N537);
nand NAND2_164 (N581, N459, N537);
nand NAND2_165 (N582, N462, N540);
nand NAND2_166 (N583, N465, N540);
nand NAND2_167 (N584, N468, N543);
nand NAND2_168 (N585, N471, N543);
nand NAND2_169 (N586, N474, N546);
nand NAND2_170 (N587, N477, N546);
nand NAND2_171 (N588, N480, N549);
nand NAND2_172 (N589, N483, N549);
nand NAND2_173 (N590, N486, N552);
nand NAND2_174 (N591, N489, N552);
nand NAND2_175 (N592, N492, N555);
nand NAND2_176 (N593, N495, N555);
nand NAND2_177 (N594, N498, N558);
nand NAND2_178 (N595, N501, N558);
nand NAND2_179 (N596, N504, N561);
nand NAND2_180 (N597, N507, N561);
nand NAND2_181 (N598, N510, N564);
nand NAND2_182 (N599, N513, N564);
nand NAND2_183 (N600, N516, N567);
nand NAND2_184 (N601, N519, N567);
nand NAND2_185 (N602, N570, N571);
nand NAND2_186 (N607, N572, N573);
nand NAND2_187 (N612, N574, N575);
nand NAND2_188 (N617, N576, N577);
nand NAND2_189 (N622, N578, N579);
nand NAND2_190 (N627, N580, N581);
nand NAND2_191 (N632, N582, N583);
nand NAND2_192 (N637, N584, N585);
nand NAND2_193 (N642, N586, N587);
nand NAND2_194 (N645, N588, N589);
nand NAND2_195 (N648, N590, N591);
nand NAND2_196 (N651, N592, N593);
nand NAND2_197 (N654, N594, N595);
nand NAND2_198 (N657, N596, N597);
nand NAND2_199 (N660, N598, N599);
nand NAND2_200 (N663, N600, N601);
nand NAND2_201 (N666, N602, N607);
nand NAND2_202 (N669, N612, N617);
nand NAND2_203 (N672, N602, N612);
nand NAND2_204 (N675, N607, N617);
nand NAND2_205 (N678, N622, N627);
nand NAND2_206 (N681, N632, N637);
nand NAND2_207 (N684, N622, N632);
nand NAND2_208 (N687, N627, N637);
nand NAND2_209 (N690, N602, N666);
nand NAND2_210 (N691, N607, N666);
nand NAND2_211 (N692, N612, N669);
nand NAND2_212 (N693, N617, N669);
nand NAND2_213 (N694, N602, N672);
nand NAND2_214 (N695, N612, N672);
nand NAND2_215 (N696, N607, N675);
nand NAND2_216 (N697, N617, N675);
nand NAND2_217 (N698, N622, N678);
nand NAND2_218 (N699, N627, N678);
nand NAND2_219 (N700, N632, N681);
nand NAND2_220 (N701, N637, N681);
nand NAND2_221 (N702, N622, N684);
nand NAND2_222 (N703, N632, N684);
nand NAND2_223 (N704, N627, N687);
nand NAND2_224 (N705, N637, N687);
nand NAND2_225 (N706, N690, N691);
nand NAND2_226 (N709, N692, N693);
nand NAND2_227 (N712, N694, N695);
nand NAND2_228 (N715, N696, N697);
nand NAND2_229 (N718, N698, N699);
nand NAND2_230 (N721, N700, N701);
nand NAND2_231 (N724, N702, N703);
nand NAND2_232 (N727, N704, N705);
nand NAND2_233 (N730, N242, N718);
nand NAND2_234 (N733, N245, N721);
nand NAND2_235 (N736, N248, N724);
nand NAND2_236 (N739, N251, N727);
nand NAND2_237 (N742, N254, N706);
nand NAND2_238 (N745, N257, N709);
nand NAND2_239 (N748, N260, N712);
nand NAND2_240 (N751, N263, N715);
nand NAND2_241 (N754, N242, N730);
nand NAND2_242 (N755, N718, N730);
nand NAND2_243 (N756, N245, N733);
nand NAND2_244 (N757, N721, N733);
nand NAND2_245 (N758, N248, N736);
nand NAND2_246 (N759, N724, N736);
nand NAND2_247 (N760, N251, N739);
nand NAND2_248 (N761, N727, N739);
nand NAND2_249 (N762, N254, N742);
nand NAND2_250 (N763, N706, N742);
nand NAND2_251 (N764, N257, N745);
nand NAND2_252 (N765, N709, N745);
nand NAND2_253 (N766, N260, N748);
nand NAND2_254 (N767, N712, N748);
nand NAND2_255 (N768, N263, N751);
nand NAND2_256 (N769, N715, N751);
nand NAND2_257 (N770, N754, N755);
nand NAND2_258 (N773, N756, N757);
nand NAND2_259 (N776, N758, N759);
nand NAND2_260 (N779, N760, N761);
nand NAND2_261 (N782, N762, N763);
nand NAND2_262 (N785, N764, N765);
nand NAND2_263 (N788, N766, N767);
nand NAND2_264 (N791, N768, N769);
nand NAND2_265 (N794, N642, N770);
nand NAND2_266 (N797, N645, N773);
nand NAND2_267 (N800, N648, N776);
nand NAND2_268 (N803, N651, N779);
nand NAND2_269 (N806, N654, N782);
nand NAND2_270 (N809, N657, N785);
nand NAND2_271 (N812, N660, N788);
nand NAND2_272 (N815, N663, N791);
nand NAND2_273 (N818, N642, N794);
nand NAND2_274 (N819, N770, N794);
nand NAND2_275 (N820, N645, N797);
nand NAND2_276 (N821, N773, N797);
nand NAND2_277 (N822, N648, N800);
nand NAND2_278 (N823, N776, N800);
nand NAND2_279 (N824, N651, N803);
nand NAND2_280 (N825, N779, N803);
nand NAND2_281 (N826, N654, N806);
nand NAND2_282 (N827, N782, N806);
nand NAND2_283 (N828, N657, N809);
nand NAND2_284 (N829, N785, N809);
nand NAND2_285 (N830, N660, N812);
nand NAND2_286 (N831, N788, N812);
nand NAND2_287 (N832, N663, N815);
nand NAND2_288 (N833, N791, N815);
nand NAND2_289 (N834, N818, N819);
nand NAND2_290 (N847, N820, N821);
nand NAND2_291 (N860, N822, N823);
nand NAND2_292 (N873, N824, N825);
nand NAND2_293 (N886, N828, N829);
nand NAND2_294 (N899, N832, N833);
nand NAND2_295 (N912, N830, N831);
nand NAND2_296 (N925, N826, N827);
not NOT1_297 (N938, N834);
not NOT1_298 (N939, N847);
not NOT1_299 (N940, N860);
not NOT1_300 (N941, N834);
not NOT1_301 (N942, N847);
not NOT1_302 (N943, N873);
not NOT1_303 (N944, N834);
not NOT1_304 (N945, N860);
not NOT1_305 (N946, N873);
not NOT1_306 (N947, N847);
not NOT1_307 (N948, N860);
not NOT1_308 (N949, N873);
not NOT1_309 (N950, N886);
not NOT1_310 (N951, N899);
not NOT1_311 (N952, N886);
not NOT1_312 (N953, N912);
not NOT1_313 (N954, N925);
not NOT1_314 (N955, N899);
not NOT1_315 (N956, N925);
not NOT1_316 (N957, N912);
not NOT1_317 (N958, N925);
not NOT1_318 (N959, N886);
not NOT1_319 (N960, N912);
not NOT1_320 (N961, N925);
not NOT1_321 (N962, N886);
not NOT1_322 (N963, N899);
not NOT1_323 (N964, N925);
not NOT1_324 (N965, N912);
not NOT1_325 (N966, N899);
not NOT1_326 (N967, N886);
not NOT1_327 (N968, N912);
not NOT1_328 (N969, N899);
not NOT1_329 (N970, N847);
not NOT1_330 (N971, N873);
not NOT1_331 (N972, N847);
not NOT1_332 (N973, N860);
not NOT1_333 (N974, N834);
not NOT1_334 (N975, N873);
not NOT1_335 (N976, N834);
not NOT1_336 (N977, N860);
and AND4_337 (N978, N938, N939, N940, N873);
and AND4_338 (N979, N941, N942, N860, N943);
and AND4_339 (N980, N944, N847, N945, N946);
and AND4_340 (N981, N834, N947, N948, N949);
and AND4_341 (N982, N958, N959, N960, N899);
and AND4_342 (N983, N961, N962, N912, N963);
and AND4_343 (N984, N964, N886, N965, N966);
and AND4_344 (N985, N925, N967, N968, N969);
or OR4_345 (N986, N978, N979, N980, N981);
or OR4_346 (N991, N982, N983, N984, N985);
and AND5_347 (N996, N925, N950, N912, N951, N986);
and AND5_348 (N1001, N925, N952, N953, N899, N986);
and AND5_349 (N1006, N954, N886, N912, N955, N986);
and AND5_350 (N1011, N956, N886, N957, N899, N986);
and AND5_351 (N1016, N834, N970, N860, N971, N991);
and AND5_352 (N1021, N834, N972, N973, N873, N991);
and AND5_353 (N1026, N974, N847, N860, N975, N991);
and AND5_354 (N1031, N976, N847, N977, N873, N991);
and AND2_355 (N1036, N834, N996);
and AND2_356 (N1039, N847, N996);
and AND2_357 (N1042, N860, N996);
and AND2_358 (N1045, N873, N996);
and AND2_359 (N1048, N834, N1001);
and AND2_360 (N1051, N847, N1001);
and AND2_361 (N1054, N860, N1001);
and AND2_362 (N1057, N873, N1001);
and AND2_363 (N1060, N834, N1006);
and AND2_364 (N1063, N847, N1006);
and AND2_365 (N1066, N860, N1006);
and AND2_366 (N1069, N873, N1006);
and AND2_367 (N1072, N834, N1011);
and AND2_368 (N1075, N847, N1011);
and AND2_369 (N1078, N860, N1011);
and AND2_370 (N1081, N873, N1011);
and AND2_371 (N1084, N925, N1016);
and AND2_372 (N1087, N886, N1016);
and AND2_373 (N1090, N912, N1016);
and AND2_374 (N1093, N899, N1016);
and AND2_375 (N1096, N925, N1021);
and AND2_376 (N1099, N886, N1021);
and AND2_377 (N1102, N912, N1021);
and AND2_378 (N1105, N899, N1021);
and AND2_379 (N1108, N925, N1026);
and AND2_380 (N1111, N886, N1026);
and AND2_381 (N1114, N912, N1026);
and AND2_382 (N1117, N899, N1026);
and AND2_383 (N1120, N925, N1031);
and AND2_384 (N1123, N886, N1031);
and AND2_385 (N1126, N912, N1031);
and AND2_386 (N1129, N899, N1031);
nand NAND2_387 (N1132, N1, N1036);
nand NAND2_388 (N1135, N8, N1039);
nand NAND2_389 (N1138, N15, N1042);
nand NAND2_390 (N1141, N22, N1045);
nand NAND2_391 (N1144, N29, N1048);
nand NAND2_392 (N1147, N36, N1051);
nand NAND2_393 (N1150, N43, N1054);
nand NAND2_394 (N1153, N50, N1057);
nand NAND2_395 (N1156, N57, N1060);
nand NAND2_396 (N1159, N64, N1063);
nand NAND2_397 (N1162, N71, N1066);
nand NAND2_398 (N1165, N78, N1069);
nand NAND2_399 (N1168, N85, N1072);
nand NAND2_400 (N1171, N92, N1075);
nand NAND2_401 (N1174, N99, N1078);
nand NAND2_402 (N1177, N106, N1081);
nand NAND2_403 (N1180, N113, N1084);
nand NAND2_404 (N1183, N120, N1087);
nand NAND2_405 (N1186, N127, N1090);
nand NAND2_406 (N1189, N134, N1093);
nand NAND2_407 (N1192, N141, N1096);
nand NAND2_408 (N1195, N148, N1099);
nand NAND2_409 (N1198, N155, N1102);
nand NAND2_410 (N1201, N162, N1105);
nand NAND2_411 (N1204, N169, N1108);
nand NAND2_412 (N1207, N176, N1111);
nand NAND2_413 (N1210, N183, N1114);
nand NAND2_414 (N1213, N190, N1117);
nand NAND2_415 (N1216, N197, N1120);
nand NAND2_416 (N1219, N204, N1123);
nand NAND2_417 (N1222, N211, N1126);
nand NAND2_418 (N1225, N218, N1129);
nand NAND2_419 (N1228, N1, N1132);
nand NAND2_420 (N1229, N1036, N1132);
nand NAND2_421 (N1230, N8, N1135);
nand NAND2_422 (N1231, N1039, N1135);
nand NAND2_423 (N1232, N15, N1138);
nand NAND2_424 (N1233, N1042, N1138);
nand NAND2_425 (N1234, N22, N1141);
nand NAND2_426 (N1235, N1045, N1141);
nand NAND2_427 (N1236, N29, N1144);
nand NAND2_428 (N1237, N1048, N1144);
nand NAND2_429 (N1238, N36, N1147);
nand NAND2_430 (N1239, N1051, N1147);
nand NAND2_431 (N1240, N43, N1150);
nand NAND2_432 (N1241, N1054, N1150);
nand NAND2_433 (N1242, N50, N1153);
nand NAND2_434 (N1243, N1057, N1153);
nand NAND2_435 (N1244, N57, N1156);
nand NAND2_436 (N1245, N1060, N1156);
nand NAND2_437 (N1246, N64, N1159);
nand NAND2_438 (N1247, N1063, N1159);
nand NAND2_439 (N1248, N71, N1162);
nand NAND2_440 (N1249, N1066, N1162);
nand NAND2_441 (N1250, N78, N1165);
nand NAND2_442 (N1251, N1069, N1165);
nand NAND2_443 (N1252, N85, N1168);
nand NAND2_444 (N1253, N1072, N1168);
nand NAND2_445 (N1254, N92, N1171);
nand NAND2_446 (N1255, N1075, N1171);
nand NAND2_447 (N1256, N99, N1174);
nand NAND2_448 (N1257, N1078, N1174);
nand NAND2_449 (N1258, N106, N1177);
nand NAND2_450 (N1259, N1081, N1177);
nand NAND2_451 (N1260, N113, N1180);
nand NAND2_452 (N1261, N1084, N1180);
nand NAND2_453 (N1262, N120, N1183);
nand NAND2_454 (N1263, N1087, N1183);
nand NAND2_455 (N1264, N127, N1186);
nand NAND2_456 (N1265, N1090, N1186);
nand NAND2_457 (N1266, N134, N1189);
nand NAND2_458 (N1267, N1093, N1189);
nand NAND2_459 (N1268, N141, N1192);
nand NAND2_460 (N1269, N1096, N1192);
nand NAND2_461 (N1270, N148, N1195);
nand NAND2_462 (N1271, N1099, N1195);
nand NAND2_463 (N1272, N155, N1198);
nand NAND2_464 (N1273, N1102, N1198);
nand NAND2_465 (N1274, N162, N1201);
nand NAND2_466 (N1275, N1105, N1201);
nand NAND2_467 (N1276, N169, N1204);
nand NAND2_468 (N1277, N1108, N1204);
nand NAND2_469 (N1278, N176, N1207);
nand NAND2_470 (N1279, N1111, N1207);
nand NAND2_471 (N1280, N183, N1210);
nand NAND2_472 (N1281, N1114, N1210);
nand NAND2_473 (N1282, N190, N1213);
nand NAND2_474 (N1283, N1117, N1213);
nand NAND2_475 (N1284, N197, N1216);
nand NAND2_476 (N1285, N1120, N1216);
nand NAND2_477 (N1286, N204, N1219);
nand NAND2_478 (N1287, N1123, N1219);
nand NAND2_479 (N1288, N211, N1222);
nand NAND2_480 (N1289, N1126, N1222);
nand NAND2_481 (N1290, N218, N1225);
nand NAND2_482 (N1291, N1129, N1225);
nand NAND2_483 (N1292, N1228, N1229);
nand NAND2_484 (N1293, N1230, N1231);
nand NAND2_485 (N1294, N1232, N1233);
nand NAND2_486 (N1295, N1234, N1235);
nand NAND2_487 (N1296, N1236, N1237);
nand NAND2_488 (N1297, N1238, N1239);
nand NAND2_489 (N1298, N1240, N1241);
nand NAND2_490 (N1299, N1242, N1243);
nand NAND2_491 (N1300, N1244, N1245);
nand NAND2_492 (N1301, N1246, N1247);
nand NAND2_493 (N1302, N1248, N1249);
nand NAND2_494 (N1303, N1250, N1251);
nand NAND2_495 (N1304, N1252, N1253);
nand NAND2_496 (N1305, N1254, N1255);
nand NAND2_497 (N1306, N1256, N1257);
nand NAND2_498 (N1307, N1258, N1259);
nand NAND2_499 (N1308, N1260, N1261);
nand NAND2_500 (N1309, N1262, N1263);
nand NAND2_501 (N1310, N1264, N1265);
nand NAND2_502 (N1311, N1266, N1267);
nand NAND2_503 (N1312, N1268, N1269);
nand NAND2_504 (N1313, N1270, N1271);
nand NAND2_505 (N1314, N1272, N1273);
nand NAND2_506 (N1315, N1274, N1275);
nand NAND2_507 (N1316, N1276, N1277);
nand NAND2_508 (N1317, N1278, N1279);
nand NAND2_509 (N1318, N1280, N1281);
nand NAND2_510 (N1319, N1282, N1283);
nand NAND2_511 (N1320, N1284, N1285);
nand NAND2_512 (N1321, N1286, N1287);
nand NAND2_513 (N1322, N1288, N1289);
nand NAND2_514 (N1323, N1290, N1291);
buf BUFF1_515 (N1324, N1292);
buf BUFF1_516 (N1325, N1293);
buf BUFF1_517 (N1326, N1294);
buf BUFF1_518 (N1327, N1295);
buf BUFF1_519 (N1328, N1296);
buf BUFF1_520 (N1329, N1297);
buf BUFF1_521 (N1330, N1298);
buf BUFF1_522 (N1331, N1299);
buf BUFF1_523 (N1332, N1300);
buf BUFF1_524 (N1333, N1301);
buf BUFF1_525 (N1334, N1302);
buf BUFF1_526 (N1335, N1303);
buf BUFF1_527 (N1336, N1304);
buf BUFF1_528 (N1337, N1305);
buf BUFF1_529 (N1338, N1306);
buf BUFF1_530 (N1339, N1307);
buf BUFF1_531 (N1340, N1308);
buf BUFF1_532 (N1341, N1309);
buf BUFF1_533 (N1342, N1310);
buf BUFF1_534 (N1343, N1311);
buf BUFF1_535 (N1344, N1312);
buf BUFF1_536 (N1345, N1313);
buf BUFF1_537 (N1346, N1314);
buf BUFF1_538 (N1347, N1315);
buf BUFF1_539 (N1348, N1316);
buf BUFF1_540 (N1349, N1317);
buf BUFF1_541 (N1350, N1318);
buf BUFF1_542 (N1351, N1319);
buf BUFF1_543 (N1352, N1320);
buf BUFF1_544 (N1353, N1321);
buf BUFF1_545 (N1354, N1322);
buf BUFF1_546 (N1355, N1323);

endmodule
